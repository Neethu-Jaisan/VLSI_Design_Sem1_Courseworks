module clk_div(
    input clk,
    output reg slow_clk
);
    reg [25:0] count = 0;

    always @(posedge clk) begin
        count <= count + 1;
        slow_clk <= count[25];
    end

endmodule
